	//********************************	 DEFINE	**************************************************
	
	`define INPUT_SIZE  			16
	
	//*******************************************************************************************
	
	module LOD
	(
	din_w,
	dout_w
	);
	
	//******************************** input & output *******************************************************

	input 		[`INPUT_SIZE-1:0]						din_w;	
	output reg	[`INPUT_SIZE-1:0]  						dout_w;
	
	//********************************************************************************
	
	reg 		[`INPUT_SIZE-1:1]						not_w;
	reg 		[`INPUT_SIZE-3:0]						and_1_w;
	reg 		[`INPUT_SIZE-2:0]						and_2_w;
	integer 	i;

	//********************************************************************************
	always @(*)
		begin
			//***************************************************************************
			not_w=~din_w[`INPUT_SIZE-1:1];
			and_1_w[`INPUT_SIZE-3]=not_w[`INPUT_SIZE-1]&not_w[`INPUT_SIZE-2];
			//***************************************************************************
			for (i=`INPUT_SIZE-2;i>=2;i=i-1)
				begin
					and_1_w[i-2]=and_1_w[i-1]&not_w[i-1];
				end			
			//***************************************************************************
			dout_w[`INPUT_SIZE-1]=din_w[`INPUT_SIZE-1];
			dout_w[`INPUT_SIZE-2]=not_w[`INPUT_SIZE-1]&din_w[`INPUT_SIZE-2];
			//***************************************************************************
			for (i=`INPUT_SIZE-3;i>=0;i=i-1)
				begin
					dout_w[i]=and_1_w[i]&din_w[i];
				end	
			//***************************************************************************
		end
	
endmodule
